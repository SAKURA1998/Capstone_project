library verilog;
use verilog.vl_types.all;
entity test1 is
end test1;
